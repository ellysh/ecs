../conf/a20-go-null.vh