# This is scenario for A20 step motor controller moving to null position

[31 47] 12
[31 71 13 05 14] 5
[31 71 12 05 14] 13
[31 71 15 32] 13
[31 72 02] 5
[31 72 02] 41
[31 44 00] 13
[31 72 01] 5
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 4
[31 72 02] 13
[31 72 02] 4
[31 72 02] 13
[31 72 02] 4
[31 72 02] 13
[31 72 02] 4
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 14
[31 72 02] 3
[31 72 02] 9
[31 72 02] 3
[31 72 02] 11
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 12
[31 72 02] 6
[31 72 02] 12
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 13
[31 72 02] 5
[31 72 02] 41
[31 42 FF FF F8 E4] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 6
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 12
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 13
[31 72 01] 5
[31 72 01] 41
[31 71 13 05 14] 13
[31 71 21 00 00 00 00] 6
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 12
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 14
[31 71 13 03 84] 3
[31 72 21] 7
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 3
[31 72 21] 10
[31 72 21] 2
[31 72 21] 12
[31 72 21] 6
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 14
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 5
[31 71 13 03 84] 12
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 6
[31 71 13 03 84] 11
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 5
[31 71 13 03 84] 13
[31 72 21] 14
[31 71 13 03 84] 3
[31 72 21] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 3
[31 72 21] 10
[31 72 21] 2
[31 72 21] 12
[31 72 21] 6
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 14
[31 71 13 03 84] 3
[31 72 21] 5
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 3
[31 72 21] 5
[31 71 13 03 84] 14
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 3
[31 72 21] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 5
[31 71 13 03 84] 7
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 14
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 14
[31 71 13 03 84] 3
[31 72 21] 5
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 14
[31 72 21] 13
[31 71 13 03 84] 3
[31 72 21] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 4
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 3
[31 72 21] 10
[31 72 21] 3
[31 72 21] 10
[31 72 21] 2
[31 72 21] 12
[31 72 21] 6
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 5
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 5
[31 71 13 03 84] 7
[31 71 13 03 84] 12
[31 72 21] 13
[31 71 13 03 84] 6
[31 72 21] 5
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 14
[31 71 13 03 84] 3
[31 72 21] 6
[31 71 13 03 84] 13
[31 72 21] 12
[31 71 13 03 84] 5
[31 72 21] 6
[31 71 13 03 84] 6
[31 71 13 03 84] 13
[31 72 21] 0
