# This is scenario to test A20 step motor controller

[31 47] 12
[31 71 13 01 F4] 10
[31 71 12 01 F4] 10
#[31 71 14 01] 10
[31 71 15 32] 13
[31 41 00] 2000
[31 47] 6
[31 41 80] 1000
[31 47] 6
#[31 41 00] 1000
#[31 47] 5
#[31 42 00 00 08 00] 10
#[31 71 14 FA] 10
