../conf/a20-test.vh